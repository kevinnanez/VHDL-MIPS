library ieee;
use ieee.std_logic_1164.all;
use work.components.all;

--y aca va el datapath
